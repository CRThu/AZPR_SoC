`timescale 1ns/100ps

`include "./Bus/bus_top.v"
`include "./Global/global_std_def.v"

module bus_top_tb;

    


endmodule // bus_top_tb